module comparador(a,b,s);
	input [31:0] a, b;
	output s;
endmodule
